../autogen/renderer.vhd