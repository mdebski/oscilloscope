../autogen/palette.vhd